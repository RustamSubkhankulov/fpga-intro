module dfa();



endmodule